// v -b js -sourcemap main.v -o hello.js

module main

fn main() {
	// Yeah... I just unlocked memories why I do not judge JavaScript for being shit

	subject := subject_create('osiris')
	username := subject.get_username()

	print('${username}')
}
